module processor;
    core core_0 (
        .clk(),

        .instr_addr(),
        .instr_in(),

        .data_we(),
        .data_addr(),
        .data_out(),
        .data_in()
    );
endmodule