module execute_unit #(
    parameter XLEN = 32,
) (

);

endmodule