typedef enum logic { alu, branch } execute_function_e;