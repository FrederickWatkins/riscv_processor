module expander (
    input [15:0] comp_instruction,

    output [31:0] exp_instruction
);
    // TODO implement decompression
endmodule
